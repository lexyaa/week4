
`timescale 1ns/1ns

module p1;

wire           clk_gen     ;

reg    [31:0]  num         ;
reg            clk         ;
reg            rst_n       ;

parameter      tCK = 1000/50;    //50MHz Clock

initial        clk = 1'b0  ;
always         #(tCK/2)
               clk = ~clk  ;

nco    dut(    .clk_gen    ( clk_gen      ),
               .num        ( 32'd50000000 ),
               .clk        ( clk          ),
               .rst_n      ( rst_n        ));

initial begin
    #(00*tCK)  rst_n = 1'b0;
    #(10*tCK)  rst_n = 1'b1;
    #(100000000*tCK)
               $finish;
end

endmodule
